class write_b_read_a_seq extends memory_virtual_sequence;
    `uvm_object_utils(write_b_read_a_seq)

    function new(string name = "write_b_read_a_seq");
        super.new(name);
    endfunction : new

    virtual task pre_start();
        super.pre_start();
        mem_sequence_b = write_seq::type_id::create("write_seq_b");
        mem_sequence_a = read_seq::type_id::create("read_seq_a");
        mem_sequence_a.same_address = 1;
    endtask : pre_start

    virtual task body();
        repeat (num) begin
            mem_sequence_b.start(p_sequencer.mem_sequencer_b);
            `uvm_info("write_b_read_a_seq", $sformatf("Writing to address: %0h", mem_sequence_b.current_addr), UVM_HIGH)
            mem_sequence_a.current_addr = mem_sequence_b.current_addr;
            mem_sequence_a.start(p_sequencer.mem_sequencer_a);
            `uvm_info("write_b_read_a_seq", $sformatf("Reading from address: %0h", mem_sequence_a.current_addr), UVM_HIGH)
        end
    endtask : body
endclass : write_b_read_a_seq