// No need to modify the memory configuration